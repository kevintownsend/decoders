module variable_length_decoder(clk, rst, push, full, size, pop, d, q);
endmodule
